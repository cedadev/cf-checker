netcdf cl_Amon_INM-CM5-0_historical_r1i1p1f1_gr1_203001-203002 {
dimensions:
        time = UNLIMITED ; // (2 currently)
        lev = 5 ;
        lat = 3 ;
        lon = 4 ;
        bnds = 2 ;
variables:
        double time(time) ;
                time:bounds = "time_bnds" ;
                time:units = "days since 2030-1-1" ;
                time:calendar = "365_day" ;
                time:axis = "T" ;
                time:long_name = "time" ;
                time:standard_name = "time" ;
        double time_bnds(time, bnds) ;
        double lev(lev) ;
                lev:bounds = "lev_bnds" ;
                lev:units = "1" ;
                lev:axis = "Z" ;
                lev:positive = "down" ;
                lev:long_name = "hybrid sigma pressure coordinate" ;
                lev:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
                lev:formula = "p = a*p0 + b*ps" ;
                lev:formula_terms = "p0: p0 a: a b: b ps: ps" ;
        double lev_bnds(lev, bnds) ;
                lev_bnds:formula = "p = a*p0 + b*ps" ;
                lev_bnds:standard_name = "atmosphere_hybrid_sigma_pressure_coordinate" ;
                lev_bnds:units = "1" ;
                lev_bnds:formula_terms = "p0: p0 a: a_bnds b: b_bnds ps: ps" ;
        double p0 ;
                p0:long_name = "vertical coordinate formula term: reference pressure" ;
                p0:units = "Pa" ;
        double a(lev) ;
                a:long_name = "vertical coordinate formula term: a(k)" ;
        double b(lev) ;
                b:long_name = "vertical coordinate formula term: b(k)" ;
        float ps(time, lat, lon) ;
                ps:long_name = "Surface Air Pressure" ;
                ps:units = "Pa" ;
        double a_bnds(lev, bnds) ;
                a_bnds:long_name = "vertical coordinate formula term: a(k+1/2)" ;
        double b_bnds(lev, bnds) ;
                b_bnds:long_name = "vertical coordinate formula term: b(k+1/2)" ;
        double lat(lat) ;
                lat:bounds = "lat_bnds" ;
                lat:units = "degrees_north" ;
                lat:axis = "Y" ;
                lat:long_name = "latitude" ;
                lat:standard_name = "latitude" ;
        double lat_bnds(lat, bnds) ;
        double lon(lon) ;
                lon:bounds = "lon_bnds" ;
                lon:units = "degrees_east" ;
                lon:axis = "X" ;
                lon:long_name = "Longitude" ;
                lon:standard_name = "longitude" ;
        double lon_bnds(lon, bnds) ;
        float cl(time, lev, lat, lon) ;
                cl:standard_name = "cloud_area_fraction_in_atmosphere_layer" ;
                cl:long_name = "Cloud Area Fraction" ;
                cl:comment = "Percentage cloud cover, including both large-scale and convective cloud." ;
                cl:units = "%" ;
                cl:original_name = "CLOUD" ;
                cl:cell_methods = "area: time: mean (interval: 20 minutes)" ;
                cl:cell_measures = "area: areacella" ;
                cl:history = "2019-04-12T14:28:43Z altered by CMOR: replaced missing value flag (1e+28) with standard missing value (1e+20). 2019-04-12T14:28:43Z altered by CMOR: Inverted axis: lev. 2019-04-12T14:28:43Z altered by CMOR: Inverted axis: lat." ;
                cl:missing_value = 1.e+20f ;
                cl:_FillValue = 1.e+20f ;

// global attributes:
                :Conventions = "CF-1.7 CMIP-6.2" ;
                :activity_id = "CMIP" ;
                :branch_method = "standard" ;
                :branch_time_in_child = 0. ;
                :branch_time_in_parent = 90885. ;
                :contact = "Evgeny Volodin (volodinev@gmail.com)" ;
                :creation_date = "2019-04-12T14:28:43Z" ;
                :data_specs_version = "01.00.27" ;
                :experiment = "all-forcing simulation of the recent past" ;
                :experiment_id = "historical" ;
                :external_variables = "areacella" ;
                :forcing_index = 1 ;
                :frequency = "mon" ;
                :further_info_url = "https://furtherinfo.es-doc.org/CMIP6.INM.INM-CM5-0.historical.none.r1i1p1f1" ;
                :grid = "gs2x1.5" ;
                :grid_label = "gr1" ;
                :history = "2019-04-12T14:28:43Z ;rewrote data to be consistent with CMIP for variable cl found in table Amon." ;
                :initialization_index = 1 ;
                :institution = "Institute for Numerical Mathematics, Russian Academy of Science, Moscow 119991, Russia" ;
                :institution_id = "INM" ;
                :mip_era = "CMIP6" ;
                :nominal_resolution = "100 km" ;
                :parent_activity_id = "CMIP" ;
                :parent_experiment_id = "piControl" ;
                :parent_mip_era = "CMIP6" ;
                :parent_source_id = "INM-CM5-0" ;
                :parent_time_units = "days since 1850-01-01" ;
                :parent_variant_label = "r1i1p1f1" ;
                :physics_index = 1 ;
                :product = "model-output" ;
                :realization_index = 1 ;
                :realm = "atmos" ;
                :references = "Clim. Dyn., 2017, 3715-3734)\'" ;
                :run_variant = "standard" ;
                :source = "INM-CM5-0 (2016): \n",
                        "aerosol: INM-AER1\n",
                        "atmos: INM-AM5-0 (2x1.5; 180 x 120 longitude/latitude; 73 levels; top level sigma = 0.0002)\n",
                        "atmosChem: none\n",
                        "land: INM-LND1\n",
                        "landIce: none\n",
                        "ocean: INM-OM5 (North Pole shifted to 60N, 90E. 0.5x0.25; 720 x 720 longitude/latitude; 40 levels; vertical sigma coordinate)\n",
                        "ocnBgchem: none\n",
                        "seaIce: INM-ICE1" ;
                :source_id = "INM-CM5-0" ;
                :source_type = "AOGCM AER" ;
                :sub_experiment = "none" ;
                :sub_experiment_id = "none" ;
                :table_id = "Amon" ;
                :table_info = "Creation Date:(30 July 2018) MD5:fa9bc503f57fb067bf398cab2c4ba77e" ;
                :title = "INM-CM5-0 output prepared for CMIP6" ;
                :tracking_id = "hdl:21.14100/8645a6fa-b7f3-4ece-ad8e-4541cee008ea" ;
                :variable_id = "cl" ;
                :variant_label = "r1i1p1f1" ;
                :license = "CMIP6 model data produced by Lawrence Livermore PCMDI is licensed under a Creative Commons Attribution ShareAlike 4.0 International License (https://creativecommons.org/licenses). Consult https://pcmdi.llnl.gov/CMIP6/TermsOfUse for terms of use governing CMIP6 output, including citation requirements and proper acknowledgment. Further information about this data, including some limitations, can be found via the further_info_url (recorded as a global attribute in this file) and at https:///pcmdi.llnl.gov/. The data producers and data providers make no warranty, either express or implied, including, but not limited to, warranties of merchantability and fitness for a particular purpose. All liabilities arising from the supply of the information (including any liability arising in negligence) are excluded to the fullest extent permitted by law." ;
                :cmor_version = "3.3.2" ;
data:

 time = 15, 45 ;

 time_bnds =
  0, 30,
  30, 60 ;

 lev = 0.899999976158142, 0.699999988079071, 0.550000011920929, 
    0.300000011920929, 0.100000001490116 ;

 lev_bnds =
  1, 0.800000011920929,
  0.800000011920929, 0.620000004768372,
  0.620000004768372, 0.419999986886978,
  0.419999986886978, 0.200000002980232,
  0.200000002980232, 0 ;

 p0 = 100000 ;

 a = 0.100000001490116, 0.219999998807907, 0.300000011920929, 
    0.200000002980232, 0.100000001490116 ;

 b = 0.800000011920929, 0.5, 0.200000002980232, 0.100000001490116, 0 ;

 ps =
  94100, 94500, 94900, 95300,
  95700, 96100, 96500, 96900,
  97300, 97700, 98100, 98500,
  94200, 94600, 95000, 95400,
  95800, 96200, 96600, 97000,
  97400, 97800, 98200, 98600 ;

 a_bnds =
  0, 0.159999996423721,
  0.159999996423721, 0.25,
  0.25, 0.25,
  0.25, 0.150000005960464,
  0.150000005960464, 0 ;

 b_bnds =
  1, 0.649999976158142,
  0.649999976158142, 0.349999994039536,
  0.349999994039536, 0.150000005960464,
  0.150000005960464, 0.0500000007450581,
  0.0500000007450581, 0 ;

 lat = 10, 20, 30 ;

 lat_bnds =
  5, 15,
  15, 25,
  25, 35 ;

 lon = 0, 90, 180, 270 ;

 lon_bnds =
  -45, 45,
  45, 135,
  135, 225,
  225, 315 ;

 cl =
  25.78, 25.86, 25.94, 26.02,
  25.46, 25.54, 25.62, 25.7,
  25.14, 25.22, 25.3, 25.38,
  24.5, 24.58, 24.66, 24.74,
  24.18, 24.26, 24.34, 24.42,
  23.86, 23.94, 24.02, 24.1,
  23.22, 23.3, 23.38, 23.46,
  22.9, 22.98, 23.06, 23.14,
  22.58, 22.66, 22.74, 22.82,
  21.94, 22.02, 22.1, 22.18,
  21.62, 21.7, 21.78, 21.86,
  21.3, 21.38, 21.46, 21.54,
  20.66, 20.74, 20.82, 20.9,
  20.34, 20.42, 20.5, 20.58,
  20.02, 20.1, 20.18, 20.26,
  25.8, 25.88, 25.96, 26.04,
  25.48, 25.56, 25.64, 25.72,
  25.16, 25.24, 25.32, 25.4,
  24.52, 24.6, 24.68, 24.76,
  24.2, 24.28, 24.36, 24.44,
  23.88, 23.96, 24.04, 24.12,
  23.24, 23.32, 23.4, 23.48,
  22.92, 23, 23.08, 23.16,
  22.6, 22.68, 22.76, 22.84,
  21.96, 22.04, 22.12, 22.2,
  21.64, 21.72, 21.8, 21.88,
  21.32, 21.4, 21.48, 21.56,
  20.68, 20.76, 20.84, 20.92,
  20.36, 20.44, 20.52, 20.6,
  20.04, 20.12, 20.2, 20.28 ;
}

